module top(	
   input wire a,
   input wire b,
   //input wire s,
   output wire f
);
   assign f=a&b;
endmodule

